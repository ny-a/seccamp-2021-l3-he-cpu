module CapitalizeString(
  input wire [255:0] my_string,
  output wire [255:0] out
);
  wire [7:0] my_string_unflattened[32];
  assign my_string_unflattened[0] = my_string[7:0];
  assign my_string_unflattened[1] = my_string[15:8];
  assign my_string_unflattened[2] = my_string[23:16];
  assign my_string_unflattened[3] = my_string[31:24];
  assign my_string_unflattened[4] = my_string[39:32];
  assign my_string_unflattened[5] = my_string[47:40];
  assign my_string_unflattened[6] = my_string[55:48];
  assign my_string_unflattened[7] = my_string[63:56];
  assign my_string_unflattened[8] = my_string[71:64];
  assign my_string_unflattened[9] = my_string[79:72];
  assign my_string_unflattened[10] = my_string[87:80];
  assign my_string_unflattened[11] = my_string[95:88];
  assign my_string_unflattened[12] = my_string[103:96];
  assign my_string_unflattened[13] = my_string[111:104];
  assign my_string_unflattened[14] = my_string[119:112];
  assign my_string_unflattened[15] = my_string[127:120];
  assign my_string_unflattened[16] = my_string[135:128];
  assign my_string_unflattened[17] = my_string[143:136];
  assign my_string_unflattened[18] = my_string[151:144];
  assign my_string_unflattened[19] = my_string[159:152];
  assign my_string_unflattened[20] = my_string[167:160];
  assign my_string_unflattened[21] = my_string[175:168];
  assign my_string_unflattened[22] = my_string[183:176];
  assign my_string_unflattened[23] = my_string[191:184];
  assign my_string_unflattened[24] = my_string[199:192];
  assign my_string_unflattened[25] = my_string[207:200];
  assign my_string_unflattened[26] = my_string[215:208];
  assign my_string_unflattened[27] = my_string[223:216];
  assign my_string_unflattened[28] = my_string[231:224];
  assign my_string_unflattened[29] = my_string[239:232];
  assign my_string_unflattened[30] = my_string[247:240];
  assign my_string_unflattened[31] = my_string[255:248];
  wire [7:0] array_index_3823;
  wire [7:0] array_index_3824;
  wire [7:0] array_index_3825;
  wire [7:0] array_index_3826;
  wire [7:0] array_index_3827;
  wire [7:0] array_index_3828;
  wire [7:0] array_index_3829;
  wire [7:0] array_index_3830;
  wire [7:0] array_index_3831;
  wire [7:0] array_index_3832;
  wire [7:0] array_index_3833;
  wire [7:0] array_index_3834;
  wire [7:0] array_index_3835;
  wire [7:0] array_index_3836;
  wire [7:0] array_index_3837;
  wire [7:0] array_index_3838;
  wire [7:0] array_index_3839;
  wire [7:0] array_index_3840;
  wire [7:0] array_index_3841;
  wire [7:0] array_index_3842;
  wire [7:0] array_index_3843;
  wire [7:0] array_index_3844;
  wire [7:0] array_index_3845;
  wire [7:0] array_index_3846;
  wire [7:0] array_index_3847;
  wire [7:0] array_index_3848;
  wire [7:0] array_index_3849;
  wire [7:0] array_index_3850;
  wire [7:0] array_index_3851;
  wire [7:0] array_index_3852;
  wire [7:0] array_index_3853;
  wire [7:0] array_index_3854;
  wire [31:0] sign_ext_3855;
  wire [31:0] sign_ext_3861;
  wire [31:0] sign_ext_3867;
  wire [31:0] sign_ext_3873;
  wire [31:0] sign_ext_3879;
  wire [31:0] sign_ext_3885;
  wire [31:0] sign_ext_3891;
  wire [31:0] sign_ext_3897;
  wire [31:0] sign_ext_3903;
  wire [31:0] sign_ext_3909;
  wire [31:0] sign_ext_3915;
  wire [31:0] sign_ext_3921;
  wire [31:0] sign_ext_3927;
  wire [31:0] sign_ext_3933;
  wire [31:0] sign_ext_3939;
  wire [31:0] sign_ext_3945;
  wire [31:0] sign_ext_3951;
  wire [31:0] sign_ext_3957;
  wire [31:0] sign_ext_3963;
  wire [31:0] sign_ext_3969;
  wire [31:0] sign_ext_3975;
  wire [31:0] sign_ext_3981;
  wire [31:0] sign_ext_3987;
  wire [31:0] sign_ext_3993;
  wire [31:0] sign_ext_3999;
  wire [31:0] sign_ext_4005;
  wire [31:0] sign_ext_4011;
  wire [31:0] sign_ext_4017;
  wire [31:0] sign_ext_4023;
  wire [31:0] sign_ext_4029;
  wire [31:0] sign_ext_4035;
  wire [31:0] sign_ext_4041;
  wire [2:0] add_4048;
  wire [2:0] add_4053;
  wire [2:0] add_4058;
  wire [2:0] add_4063;
  wire [2:0] add_4068;
  wire [2:0] add_4073;
  wire [2:0] add_4078;
  wire [2:0] add_4083;
  wire [2:0] add_4088;
  wire [2:0] add_4093;
  wire [2:0] add_4098;
  wire [2:0] add_4103;
  wire [2:0] add_4108;
  wire [2:0] add_4113;
  wire [2:0] add_4118;
  wire [2:0] add_4123;
  wire [2:0] add_4128;
  wire [2:0] add_4133;
  wire [2:0] add_4138;
  wire [2:0] add_4143;
  wire [2:0] add_4148;
  wire [2:0] add_4153;
  wire [2:0] add_4158;
  wire [2:0] add_4163;
  wire [2:0] add_4168;
  wire [2:0] add_4173;
  wire [2:0] add_4178;
  wire [2:0] add_4183;
  wire [2:0] add_4188;
  wire [2:0] add_4193;
  wire [2:0] add_4198;
  wire [2:0] add_4203;
  wire [7:0] array_4301[32];
  assign array_index_3823 = my_string_unflattened[32'h0000_0000];
  assign array_index_3824 = my_string_unflattened[32'h0000_0001];
  assign array_index_3825 = my_string_unflattened[32'h0000_0002];
  assign array_index_3826 = my_string_unflattened[32'h0000_0003];
  assign array_index_3827 = my_string_unflattened[32'h0000_0004];
  assign array_index_3828 = my_string_unflattened[32'h0000_0005];
  assign array_index_3829 = my_string_unflattened[32'h0000_0006];
  assign array_index_3830 = my_string_unflattened[32'h0000_0007];
  assign array_index_3831 = my_string_unflattened[32'h0000_0008];
  assign array_index_3832 = my_string_unflattened[32'h0000_0009];
  assign array_index_3833 = my_string_unflattened[32'h0000_000a];
  assign array_index_3834 = my_string_unflattened[32'h0000_000b];
  assign array_index_3835 = my_string_unflattened[32'h0000_000c];
  assign array_index_3836 = my_string_unflattened[32'h0000_000d];
  assign array_index_3837 = my_string_unflattened[32'h0000_000e];
  assign array_index_3838 = my_string_unflattened[32'h0000_000f];
  assign array_index_3839 = my_string_unflattened[32'h0000_0010];
  assign array_index_3840 = my_string_unflattened[32'h0000_0011];
  assign array_index_3841 = my_string_unflattened[32'h0000_0012];
  assign array_index_3842 = my_string_unflattened[32'h0000_0013];
  assign array_index_3843 = my_string_unflattened[32'h0000_0014];
  assign array_index_3844 = my_string_unflattened[32'h0000_0015];
  assign array_index_3845 = my_string_unflattened[32'h0000_0016];
  assign array_index_3846 = my_string_unflattened[32'h0000_0017];
  assign array_index_3847 = my_string_unflattened[32'h0000_0018];
  assign array_index_3848 = my_string_unflattened[32'h0000_0019];
  assign array_index_3849 = my_string_unflattened[32'h0000_001a];
  assign array_index_3850 = my_string_unflattened[32'h0000_001b];
  assign array_index_3851 = my_string_unflattened[32'h0000_001c];
  assign array_index_3852 = my_string_unflattened[32'h0000_001d];
  assign array_index_3853 = my_string_unflattened[32'h0000_001e];
  assign array_index_3854 = my_string_unflattened[32'h0000_001f];
  assign sign_ext_3855 = {{24{array_index_3823[7]}}, array_index_3823};
  assign sign_ext_3861 = {{24{array_index_3824[7]}}, array_index_3824};
  assign sign_ext_3867 = {{24{array_index_3825[7]}}, array_index_3825};
  assign sign_ext_3873 = {{24{array_index_3826[7]}}, array_index_3826};
  assign sign_ext_3879 = {{24{array_index_3827[7]}}, array_index_3827};
  assign sign_ext_3885 = {{24{array_index_3828[7]}}, array_index_3828};
  assign sign_ext_3891 = {{24{array_index_3829[7]}}, array_index_3829};
  assign sign_ext_3897 = {{24{array_index_3830[7]}}, array_index_3830};
  assign sign_ext_3903 = {{24{array_index_3831[7]}}, array_index_3831};
  assign sign_ext_3909 = {{24{array_index_3832[7]}}, array_index_3832};
  assign sign_ext_3915 = {{24{array_index_3833[7]}}, array_index_3833};
  assign sign_ext_3921 = {{24{array_index_3834[7]}}, array_index_3834};
  assign sign_ext_3927 = {{24{array_index_3835[7]}}, array_index_3835};
  assign sign_ext_3933 = {{24{array_index_3836[7]}}, array_index_3836};
  assign sign_ext_3939 = {{24{array_index_3837[7]}}, array_index_3837};
  assign sign_ext_3945 = {{24{array_index_3838[7]}}, array_index_3838};
  assign sign_ext_3951 = {{24{array_index_3839[7]}}, array_index_3839};
  assign sign_ext_3957 = {{24{array_index_3840[7]}}, array_index_3840};
  assign sign_ext_3963 = {{24{array_index_3841[7]}}, array_index_3841};
  assign sign_ext_3969 = {{24{array_index_3842[7]}}, array_index_3842};
  assign sign_ext_3975 = {{24{array_index_3843[7]}}, array_index_3843};
  assign sign_ext_3981 = {{24{array_index_3844[7]}}, array_index_3844};
  assign sign_ext_3987 = {{24{array_index_3845[7]}}, array_index_3845};
  assign sign_ext_3993 = {{24{array_index_3846[7]}}, array_index_3846};
  assign sign_ext_3999 = {{24{array_index_3847[7]}}, array_index_3847};
  assign sign_ext_4005 = {{24{array_index_3848[7]}}, array_index_3848};
  assign sign_ext_4011 = {{24{array_index_3849[7]}}, array_index_3849};
  assign sign_ext_4017 = {{24{array_index_3850[7]}}, array_index_3850};
  assign sign_ext_4023 = {{24{array_index_3851[7]}}, array_index_3851};
  assign sign_ext_4029 = {{24{array_index_3852[7]}}, array_index_3852};
  assign sign_ext_4035 = {{24{array_index_3853[7]}}, array_index_3853};
  assign sign_ext_4041 = {{24{array_index_3854[7]}}, array_index_3854};
  assign add_4048 = array_index_3823[7:5] + 3'h7;
  assign add_4053 = array_index_3824[7:5] + 3'h7;
  assign add_4058 = array_index_3825[7:5] + 3'h7;
  assign add_4063 = array_index_3826[7:5] + 3'h7;
  assign add_4068 = array_index_3827[7:5] + 3'h7;
  assign add_4073 = array_index_3828[7:5] + 3'h7;
  assign add_4078 = array_index_3829[7:5] + 3'h7;
  assign add_4083 = array_index_3830[7:5] + 3'h7;
  assign add_4088 = array_index_3831[7:5] + 3'h7;
  assign add_4093 = array_index_3832[7:5] + 3'h7;
  assign add_4098 = array_index_3833[7:5] + 3'h7;
  assign add_4103 = array_index_3834[7:5] + 3'h7;
  assign add_4108 = array_index_3835[7:5] + 3'h7;
  assign add_4113 = array_index_3836[7:5] + 3'h7;
  assign add_4118 = array_index_3837[7:5] + 3'h7;
  assign add_4123 = array_index_3838[7:5] + 3'h7;
  assign add_4128 = array_index_3839[7:5] + 3'h7;
  assign add_4133 = array_index_3840[7:5] + 3'h7;
  assign add_4138 = array_index_3841[7:5] + 3'h7;
  assign add_4143 = array_index_3842[7:5] + 3'h7;
  assign add_4148 = array_index_3843[7:5] + 3'h7;
  assign add_4153 = array_index_3844[7:5] + 3'h7;
  assign add_4158 = array_index_3845[7:5] + 3'h7;
  assign add_4163 = array_index_3846[7:5] + 3'h7;
  assign add_4168 = array_index_3847[7:5] + 3'h7;
  assign add_4173 = array_index_3848[7:5] + 3'h7;
  assign add_4178 = array_index_3849[7:5] + 3'h7;
  assign add_4183 = array_index_3850[7:5] + 3'h7;
  assign add_4188 = array_index_3851[7:5] + 3'h7;
  assign add_4193 = array_index_3852[7:5] + 3'h7;
  assign add_4198 = array_index_3853[7:5] + 3'h7;
  assign add_4203 = array_index_3854[7:5] + 3'h7;
  assign array_4301[0] = ($signed(sign_ext_3855) >= $signed(32'h0000_0061) & $signed(sign_ext_3855) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3823 : {add_4048, array_index_3823[4:0]};
  assign array_4301[1] = (sign_ext_3855 == 32'h0000_0020 & $signed(sign_ext_3861) >= $signed(32'h0000_0061) & $signed(sign_ext_3861) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3824 : {add_4053, array_index_3824[4:0]};
  assign array_4301[2] = (sign_ext_3861 == 32'h0000_0020 & $signed(sign_ext_3867) >= $signed(32'h0000_0061) & $signed(sign_ext_3867) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3825 : {add_4058, array_index_3825[4:0]};
  assign array_4301[3] = (sign_ext_3867 == 32'h0000_0020 & $signed(sign_ext_3873) >= $signed(32'h0000_0061) & $signed(sign_ext_3873) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3826 : {add_4063, array_index_3826[4:0]};
  assign array_4301[4] = (sign_ext_3873 == 32'h0000_0020 & $signed(sign_ext_3879) >= $signed(32'h0000_0061) & $signed(sign_ext_3879) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3827 : {add_4068, array_index_3827[4:0]};
  assign array_4301[5] = (sign_ext_3879 == 32'h0000_0020 & $signed(sign_ext_3885) >= $signed(32'h0000_0061) & $signed(sign_ext_3885) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3828 : {add_4073, array_index_3828[4:0]};
  assign array_4301[6] = (sign_ext_3885 == 32'h0000_0020 & $signed(sign_ext_3891) >= $signed(32'h0000_0061) & $signed(sign_ext_3891) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3829 : {add_4078, array_index_3829[4:0]};
  assign array_4301[7] = (sign_ext_3891 == 32'h0000_0020 & $signed(sign_ext_3897) >= $signed(32'h0000_0061) & $signed(sign_ext_3897) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3830 : {add_4083, array_index_3830[4:0]};
  assign array_4301[8] = (sign_ext_3897 == 32'h0000_0020 & $signed(sign_ext_3903) >= $signed(32'h0000_0061) & $signed(sign_ext_3903) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3831 : {add_4088, array_index_3831[4:0]};
  assign array_4301[9] = (sign_ext_3903 == 32'h0000_0020 & $signed(sign_ext_3909) >= $signed(32'h0000_0061) & $signed(sign_ext_3909) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3832 : {add_4093, array_index_3832[4:0]};
  assign array_4301[10] = (sign_ext_3909 == 32'h0000_0020 & $signed(sign_ext_3915) >= $signed(32'h0000_0061) & $signed(sign_ext_3915) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3833 : {add_4098, array_index_3833[4:0]};
  assign array_4301[11] = (sign_ext_3915 == 32'h0000_0020 & $signed(sign_ext_3921) >= $signed(32'h0000_0061) & $signed(sign_ext_3921) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3834 : {add_4103, array_index_3834[4:0]};
  assign array_4301[12] = (sign_ext_3921 == 32'h0000_0020 & $signed(sign_ext_3927) >= $signed(32'h0000_0061) & $signed(sign_ext_3927) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3835 : {add_4108, array_index_3835[4:0]};
  assign array_4301[13] = (sign_ext_3927 == 32'h0000_0020 & $signed(sign_ext_3933) >= $signed(32'h0000_0061) & $signed(sign_ext_3933) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3836 : {add_4113, array_index_3836[4:0]};
  assign array_4301[14] = (sign_ext_3933 == 32'h0000_0020 & $signed(sign_ext_3939) >= $signed(32'h0000_0061) & $signed(sign_ext_3939) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3837 : {add_4118, array_index_3837[4:0]};
  assign array_4301[15] = (sign_ext_3939 == 32'h0000_0020 & $signed(sign_ext_3945) >= $signed(32'h0000_0061) & $signed(sign_ext_3945) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3838 : {add_4123, array_index_3838[4:0]};
  assign array_4301[16] = (sign_ext_3945 == 32'h0000_0020 & $signed(sign_ext_3951) >= $signed(32'h0000_0061) & $signed(sign_ext_3951) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3839 : {add_4128, array_index_3839[4:0]};
  assign array_4301[17] = (sign_ext_3951 == 32'h0000_0020 & $signed(sign_ext_3957) >= $signed(32'h0000_0061) & $signed(sign_ext_3957) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3840 : {add_4133, array_index_3840[4:0]};
  assign array_4301[18] = (sign_ext_3957 == 32'h0000_0020 & $signed(sign_ext_3963) >= $signed(32'h0000_0061) & $signed(sign_ext_3963) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3841 : {add_4138, array_index_3841[4:0]};
  assign array_4301[19] = (sign_ext_3963 == 32'h0000_0020 & $signed(sign_ext_3969) >= $signed(32'h0000_0061) & $signed(sign_ext_3969) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3842 : {add_4143, array_index_3842[4:0]};
  assign array_4301[20] = (sign_ext_3969 == 32'h0000_0020 & $signed(sign_ext_3975) >= $signed(32'h0000_0061) & $signed(sign_ext_3975) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3843 : {add_4148, array_index_3843[4:0]};
  assign array_4301[21] = (sign_ext_3975 == 32'h0000_0020 & $signed(sign_ext_3981) >= $signed(32'h0000_0061) & $signed(sign_ext_3981) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3844 : {add_4153, array_index_3844[4:0]};
  assign array_4301[22] = (sign_ext_3981 == 32'h0000_0020 & $signed(sign_ext_3987) >= $signed(32'h0000_0061) & $signed(sign_ext_3987) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3845 : {add_4158, array_index_3845[4:0]};
  assign array_4301[23] = (sign_ext_3987 == 32'h0000_0020 & $signed(sign_ext_3993) >= $signed(32'h0000_0061) & $signed(sign_ext_3993) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3846 : {add_4163, array_index_3846[4:0]};
  assign array_4301[24] = (sign_ext_3993 == 32'h0000_0020 & $signed(sign_ext_3999) >= $signed(32'h0000_0061) & $signed(sign_ext_3999) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3847 : {add_4168, array_index_3847[4:0]};
  assign array_4301[25] = (sign_ext_3999 == 32'h0000_0020 & $signed(sign_ext_4005) >= $signed(32'h0000_0061) & $signed(sign_ext_4005) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3848 : {add_4173, array_index_3848[4:0]};
  assign array_4301[26] = (sign_ext_4005 == 32'h0000_0020 & $signed(sign_ext_4011) >= $signed(32'h0000_0061) & $signed(sign_ext_4011) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3849 : {add_4178, array_index_3849[4:0]};
  assign array_4301[27] = (sign_ext_4011 == 32'h0000_0020 & $signed(sign_ext_4017) >= $signed(32'h0000_0061) & $signed(sign_ext_4017) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3850 : {add_4183, array_index_3850[4:0]};
  assign array_4301[28] = (sign_ext_4017 == 32'h0000_0020 & $signed(sign_ext_4023) >= $signed(32'h0000_0061) & $signed(sign_ext_4023) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3851 : {add_4188, array_index_3851[4:0]};
  assign array_4301[29] = (sign_ext_4023 == 32'h0000_0020 & $signed(sign_ext_4029) >= $signed(32'h0000_0061) & $signed(sign_ext_4029) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3852 : {add_4193, array_index_3852[4:0]};
  assign array_4301[30] = (sign_ext_4029 == 32'h0000_0020 & $signed(sign_ext_4035) >= $signed(32'h0000_0061) & $signed(sign_ext_4035) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3853 : {add_4198, array_index_3853[4:0]};
  assign array_4301[31] = (sign_ext_4035 == 32'h0000_0020 & $signed(sign_ext_4041) >= $signed(32'h0000_0061) & $signed(sign_ext_4041) <= $signed(32'h0000_007a)) == 1'h0 ? array_index_3854 : {add_4203, array_index_3854[4:0]};
  assign out = {array_4301[31], array_4301[30], array_4301[29], array_4301[28], array_4301[27], array_4301[26], array_4301[25], array_4301[24], array_4301[23], array_4301[22], array_4301[21], array_4301[20], array_4301[19], array_4301[18], array_4301[17], array_4301[16], array_4301[15], array_4301[14], array_4301[13], array_4301[12], array_4301[11], array_4301[10], array_4301[9], array_4301[8], array_4301[7], array_4301[6], array_4301[5], array_4301[4], array_4301[3], array_4301[2], array_4301[1], array_4301[0]};
endmodule
